
`define	RA			3'b101
`define	RSUB			3'b001
`define	RADD			3'b010	
`define	RSUBMUL			6'b000
`define	RBEQ			6'b100				
`define	RMUL			3'b110
`define	RADDMUL			3'b111
`define	RBNE			6'b011
